-- Projet de stage ING4 : RISC-V
-- ECE Paris / ARESIA
-- BOOTLOADER VHDL

-- LIBRARIES
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- ENTITY
entity Bootloader is
	port (
		--INPUTS
		clk 					: in std_logic;
		CS 					: in std_logic; 							--chip select
		addrInstBoot		: in std_logic_vector(11 downto 0); --addr of boot instruction
		--OUTPUT
		instBoot				: out std_logic_vector(31 downto 0)    --output boot instruction
	);
end entity;

-- ARCHITECTURE
architecture archi of Bootloader is
--	TYPE ROM IS ARRAY(0 TO 71) OF std_logic_vector(0 to 31);
--	TYPE ROM IS ARRAY(0 TO 211) OF std_logic_vector(0 to 31);
	TYPE ROM IS ARRAY(0 TO 215) OF std_logic_vector(0 to 31);
--	TYPE ROM IS ARRAY(0 TO 214) OF std_logic_vector(0 to 31);


	SIGNAL rom_block : ROM :=(
--		x"00001137" , x"00c000ef" , x"00100073" , x"0000006f" , x"80000737" , x"000107b7" , x"fff78793" , x"00f72423",
--		x"83c0c7b7" , x"08778793" , x"00f72223" , x"01800693" , x"00000313" , x"c0000737" , x"ff800613" , x"00072783",
--		x"0047f793" , x"fe078ce3" , x"00472783" , x"00072503" , x"00157513" , x"fe051ce3" , x"00f72223" , x"00d797b3",
--		x"00f36333" , x"ff868693" , x"fcc69ae3" , x"08030263" , x"fffffe37" , x"004e0e13" , x"01c30e33" , x"00030893",
--		x"c0000737" , x"ff800813" , x"00c0006f" , x"06088263" , x"071e0063" , x"41130633" , x"00050593" , x"01800693",
--		x"00072783" , x"0047f793" , x"fe078ce3" , x"00472783" , x"00d797b3" , x"00f5e5b3" , x"ff868693" , x"ff0692e3",
--		x"ffc88893" , x"00b62023" , x"01800693" , x"00d5d633" , x"0ff67613" , x"00072783" , x"0017f793" , x"fe079ce3",
--		x"00c72223" , x"ff868693" , x"ff0692e3" , x"fa1ff06f" , x"00000693" , x"c0000737" , x"00001637" , x"ffc60613",
--		x"00072783" , x"0017f793" , x"fe079ce3" , x"0006c783" , x"00f72223" , x"00168693" , x"fec694e3" , x"0000006f"
		
		-- no wait no debug 211
--		x"00001137" , x"198000ef" , x"00100073" , x"0000006f" , x"ff010113" , x"00012623" , x"00a05e63" , x"00000713",
--		x"00c12783" , x"00178793" , x"00f12623" , x"00170713" , x"fee518e3" , x"00012623" , x"01010113" , x"00008067",
--		x"fe050513" , x"0ff57713" , x"03f00793" , x"14e7e063" , x"00271513" , x"25000793" , x"00f50533" , x"00052783",
--		x"00078067" , x"0f900513" , x"00008067" , x"0a400513" , x"00008067" , x"0b000513" , x"00008067" , x"09900513",
--		x"00008067" , x"09200513" , x"00008067" , x"08200513" , x"00008067" , x"0f800513" , x"00008067" , x"08000513",
--		x"00008067" , x"09000513" , x"00008067" , x"08800513" , x"00008067" , x"08300513" , x"00008067" , x"0c600513",
--		x"00008067" , x"0a100513" , x"00008067" , x"08600513" , x"00008067" , x"08e00513" , x"00008067" , x"0c200513",
--		x"00008067" , x"08b00513" , x"00008067" , x"0e100513" , x"00008067" , x"08a00513" , x"00008067" , x"0c700513",
--		x"00008067" , x"0aa00513" , x"00008067" , x"0ab00513" , x"00008067" , x"08c00513" , x"00008067" , x"09800513",
--		x"00008067" , x"0ce00513" , x"00008067" , x"09200513" , x"00008067" , x"08700513" , x"00008067" , x"0c100513",
--		x"00008067" , x"0b500513" , x"00008067" , x"09500513" , x"00008067" , x"08900513" , x"00008067" , x"09100513",
--		x"00008067" , x"0a400513" , x"00008067" , x"0ff00513" , x"00008067" , x"07f00513" , x"00008067" , x"0bf00513",
--		x"00008067" , x"0f700513" , x"00008067" , x"07f00513" , x"00008067" , x"0c000513" , x"00008067" , x"fd010113",
--		x"02112623" , x"02812423" , x"02912223" , x"03212023" , x"01312e23" , x"80000737" , x"000107b7" , x"fff78793",
--		x"00f72423" , x"83c0c7b7" , x"08778793" , x"00f72223" , x"444347b7" , x"24178793" , x"00f12223" , x"484747b7",
--		x"64578793" , x"00f12423" , x"4c4b57b7" , x"a4978793" , x"00f12623" , x"00414783" , x"0ff7f793" , x"04c00713",
--		x"04e78663" , x"00000413" , x"800009b7" , x"04c00913" , x"00040793" , x"00140413" , x"01040713" , x"002704b3",
--		x"ff44c703" , x"0ff77713" , x"01078793" , x"002787b3" , x"fee78a23" , x"ff47c503" , x"e09ff0ef" , x"00a9a223",
--		x"ff44c783" , x"0ff7f793" , x"fd2794e3" , x"0000006f" , x"0000016c" , x"0000018c" , x"0000018c" , x"0000018c",
--		x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c",
--		x"0000018c" , x"0000017c" , x"00000174" , x"0000018c" , x"00000194" , x"00000064" , x"0000006c" , x"00000074",
--		x"0000007c" , x"00000084" , x"0000008c" , x"00000094" , x"0000009c" , x"000000a4" , x"0000018c" , x"0000018c",
--		x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"000000ac" , x"000000b4" , x"000000bc",
--		x"000000c4" , x"000000cc" , x"000000d4" , x"000000dc" , x"000000e4" , x"00000064" , x"000000ec" , x"000000f4",
--		x"000000fc" , x"00000104" , x"0000010c" , x"00000194" , x"00000114" , x"0000011c" , x"00000124" , x"0000012c",
--		x"00000134" , x"0000013c" , x"00000144" , x"0000014c" , x"00000154" , x"0000015c" , x"00000164" , x"0000018c",
--		x"0000018c" , x"0000018c" , x"0000018c" , x"00000184"

		-- no wait with debug
		x"00001137" , x"198000ef" , x"00100073" , x"0000006f" , x"ff010113" , x"00012623" , x"00a05e63" , x"00000713",
		x"00c12783" , x"00178793" , x"00f12623" , x"00170713" , x"fee518e3" , x"00012623" , x"01010113" , x"00008067",
		x"fe050513" , x"0ff57713" , x"03f00793" , x"14e7e063" , x"00271513" , x"26000793" , x"00f50533" , x"00052783",
		x"00078067" , x"0f900513" , x"00008067" , x"0a400513" , x"00008067" , x"0b000513" , x"00008067" , x"09900513",
		x"00008067" , x"09200513" , x"00008067" , x"08200513" , x"00008067" , x"0f800513" , x"00008067" , x"08000513",
		x"00008067" , x"09000513" , x"00008067" , x"08800513" , x"00008067" , x"08300513" , x"00008067" , x"0c600513",
		x"00008067" , x"0a100513" , x"00008067" , x"08600513" , x"00008067" , x"08e00513" , x"00008067" , x"0c200513",
		x"00008067" , x"08b00513" , x"00008067" , x"0e100513" , x"00008067" , x"08a00513" , x"00008067" , x"0c700513",
		x"00008067" , x"0aa00513" , x"00008067" , x"0ab00513" , x"00008067" , x"08c00513" , x"00008067" , x"09800513",
		x"00008067" , x"0ce00513" , x"00008067" , x"09200513" , x"00008067" , x"08700513" , x"00008067" , x"0c100513",
		x"00008067" , x"0b500513" , x"00008067" , x"09500513" , x"00008067" , x"08900513" , x"00008067" , x"09100513",
		x"00008067" , x"0a400513" , x"00008067" , x"0ff00513" , x"00008067" , x"07f00513" , x"00008067" , x"0bf00513",
		x"00008067" , x"0f700513" , x"00008067" , x"07f00513" , x"00008067" , x"0c000513" , x"00008067" , x"fd010113",
		x"02112623" , x"02812423" , x"02912223" , x"03212023" , x"01312e23" , x"80000737" , x"01072783" , x"2007f793",
		x"fe078ce3" , x"80000737" , x"000107b7" , x"fff78793" , x"00f72423" , x"83c0c7b7" , x"08778793" , x"00f72223",
		x"444347b7" , x"24178793" , x"00f12223" , x"484747b7" , x"64578793" , x"00f12423" , x"4c4b57b7" , x"a4978793",
		x"00f12623" , x"00414783" , x"0ff7f793" , x"04c00713" , x"04e78663" , x"00000413" , x"800009b7" , x"04c00913",
		x"00040793" , x"00140413" , x"01040713" , x"002704b3" , x"ff44c703" , x"0ff77713" , x"01078793" , x"002787b3",
		x"fee78a23" , x"ff47c503" , x"df9ff0ef" , x"00a9a223" , x"ff44c783" , x"0ff7f793" , x"fd2794e3" , x"0000006f",
		x"0000016c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c",
		x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000017c" , x"00000174" , x"0000018c",
		x"00000194" , x"00000064" , x"0000006c" , x"00000074" , x"0000007c" , x"00000084" , x"0000008c" , x"00000094",
		x"0000009c" , x"000000a4" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c",
		x"0000018c" , x"000000ac" , x"000000b4" , x"000000bc" , x"000000c4" , x"000000cc" , x"000000d4" , x"000000dc",
		x"000000e4" , x"00000064" , x"000000ec" , x"000000f4" , x"000000fc" , x"00000104" , x"0000010c" , x"00000194",
		x"00000114" , x"0000011c" , x"00000124" , x"0000012c" , x"00000134" , x"0000013c" , x"00000144" , x"0000014c",
		x"00000154" , x"0000015c" , x"00000164" , x"0000018c" , x"0000018c" , x"0000018c" , x"0000018c" , x"00000184"
		

		
		
	);
	
	signal sigad : integer;
	signal sigpc : std_logic_vector(11 downto 0);
	
	begin
		sigpc <= addrInstBoot(11 downto 0);
		instBoot <= rom_block(sigad) when rising_edge(clk);
		sigad <= 215 when ((unsigned(sigpc) > 215)) else to_integer(unsigned(sigpc));
	
end archi;
-- END FILE